module IO_mod_robot
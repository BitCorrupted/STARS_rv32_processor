`timescale 1ms/10ps
module tb_request_unit();




endmodule